module Register1Bit 
(
			input Clk, Reset, D,
			output logic Q
);

always_ff @ (posedge Clk)
begin
	if(Reset)
		Q <= 1'b0;
	else
		Q <= D;
end
endmodule
