
module  SRAM_Controller
(
		input logic Clk,
		





);

enum logic[3:0]

always_ff @ (posedge Clk)
begin
		
end
	
	
always_comb
begin






end
	
endmodule
