
module  finalProjectTopLevel( input         CLOCK_50,
                       input[3:0]    KEY, //bit 0 is set up as Reset
							  output [6:0]  HEX0, HEX1,// HEX2, HEX3, HEX4, HEX5, HEX6, HEX7,
							  //output [8:0]  LEDG,
							  //output [17:0] LEDR,
							  // VGA Interface
                       output [7:0]  VGA_R,					//VGA Red
							                VGA_G,					//VGA Green
												 VGA_B,					//VGA Blue
							  output        VGA_CLK,				//VGA Clock
							                VGA_SYNC_N,			//VGA Sync signal
												 VGA_BLANK_N,			//VGA Blank signal
												 VGA_VS,					//VGA virtical sync signal
												 VGA_HS,					//VGA horizontal sync signal
							  // CY7C67200 Interface
							  inout [15:0]  OTG_DATA,						//	CY7C67200 Data bus 16 Bits
							  output [1:0]  OTG_ADDR,						//	CY7C67200 Address 2 Bits
							  output        OTG_CS_N,						//	CY7C67200 Chip Select
												 OTG_RD_N,						//	CY7C67200 Write
												 OTG_WR_N,						//	CY7C67200 Read
												 OTG_RST_N,						//	CY7C67200 Reset
							  input			 OTG_INT,						//	CY7C67200 Interrupt
							  // SDRAM Interface for Nios II Software
							  output [12:0] DRAM_ADDR,				// SDRAM Address 13 Bits
							  inout [31:0]  DRAM_DQ,				// SDRAM Data 32 Bits
							  output [1:0]  DRAM_BA,				// SDRAM Bank Address 2 Bits
							  output [3:0]  DRAM_DQM,				// SDRAM Data Mast 4 Bits
							  output			 DRAM_RAS_N,			// SDRAM Row Address Strobe
							  output			 DRAM_CAS_N,			// SDRAM Column Address Strobe
							  output			 DRAM_CKE,				// SDRAM Clock Enable
							  output			 DRAM_WE_N,				// SDRAM Write Enable
							  output			 DRAM_CS_N,				// SDRAM Chip Select
							  output			 DRAM_CLK				// SDRAM Clock
											);

    logic Reset_h, Reset_sh, vssig, Clk;
    logic [9:0] drawxsig, drawysig, ballxsig, ballysig, ballsizesig;
	logic [15:0] keycode;

	logic [5:0]colorValue;
	logic [15:0] colorCounter;
	logic [1:0] gameStateWire;

	assign Clk = CLOCK_50;
    assign {Reset_h}=~ (KEY[0]);  // The push buttons are active low
	assign {Reset_sh}=~ (KEY[3]);  // The push buttons are active low

	 wire [1:0] hpi_addr;
	 wire [15:0] hpi_data_in, hpi_data_out;
	 wire hpi_r, hpi_w,hpi_cs;

	 hpi_io_intf hpi_io_inst
	 (
										 .from_sw_address(hpi_addr),
										 .from_sw_data_in(hpi_data_in),
										 .from_sw_data_out(hpi_data_out),
										 .from_sw_r(hpi_r),
										 .from_sw_w(hpi_w),
										 .from_sw_cs(hpi_cs),
		 								 .OTG_DATA(OTG_DATA),
										 .OTG_ADDR(OTG_ADDR),
										 .OTG_RD_N(OTG_RD_N),
										 .OTG_WR_N(OTG_WR_N),
										 .OTG_CS_N(OTG_CS_N),
										 .OTG_RST_N(OTG_RST_N),
										 .OTG_INT(OTG_INT),
										 .Clk(Clk),
										 .Reset(Reset_h)
	 );

	 //The connections for nios_system might be named different depending on how you set up Qsys
	 nios_system nios_system
	 (
										 .clk_clk(Clk),
										 .reset_reset_n(KEY[0]),
										 .sdram_wire_addr(DRAM_ADDR),
										 .sdram_wire_ba(DRAM_BA),
										 .sdram_wire_cas_n(DRAM_CAS_N),
										 .sdram_wire_cke(DRAM_CKE),
										 .sdram_wire_cs_n(DRAM_CS_N),
										 .sdram_wire_dq(DRAM_DQ),
										 .sdram_wire_dqm(DRAM_DQM),
										 .sdram_wire_ras_n(DRAM_RAS_N),
										 .sdram_wire_we_n(DRAM_WE_N),
										 .sdram_out_clk(DRAM_CLK),
										 .keycode_export(keycode),
										 .otg_hpi_address_export(hpi_addr),
										 .otg_hpi_data_in_port(hpi_data_in),
										 .otg_hpi_data_out_port(hpi_data_out),
										 .otg_hpi_cs_export(hpi_cs),
										 .otg_hpi_r_export(hpi_r),
										 .otg_hpi_w_export(hpi_w)
	);

	//Fill in the connections for the rest of the modules
    vga_controller vgasync_instance
	 (
										.Clk(Clk),
										.Reset(Reset_sh),
										.hs(VGA_HS),
										.vs(VGA_VS),
										.pixel_clk(VGA_CLK),
										.blank(VGA_BLANK_N),
										.sync(VGA_SYNC_N),
										.DrawX(drawxsig),
										.DrawY(drawysig)

	 );


    Color_Mapper8Bit color_instance
	 (
										.Clk(Clk),
										.memMappedValue(colorValue),
										.Red(VGA_R),
										.Green(VGA_G),
										.Blue(VGA_B)
	 );

	GameController gameControllerInst
	(
										.Clk(Clk),
										.Reset(Reset_sh),
										.keycode(keycode),
										.playerDead(),
										.gameState(gameStateWire)
	);

	GameEngine	gameEngineInst
	(
                    s

	);




	/*
	SIMPLE STATE MACHINE TO TEST GAME STATE CONTROLLER

	always_ff @ (posedge Clk)
	begin
		if(gameStateWire == 2'b01)		// if we are in the play state
		begin
			if(colorValue == 6'h3C || VGA_VS == 1'b0)
				begin
					colorValue <= 6'h00;
					colorCounter <= 16'b0000;
				end
			else if(colorCounter == 16'h36B0)
				begin
					colorValue <= colorValue + 6'h01;
					colorCounter <= 16'b0000;
				end
			else
				colorCounter <= colorCounter + 16'b0001;
		end
		else
		begin
				colorValue <= 6'h00;
				colorCounter <= 16'b0000;
		end
	end
	*/

	 HexDriver hex_inst_0 (keycode[3:0], HEX0);
	 HexDriver hex_inst_1 (keycode[7:4], HEX1);


	 /**************************************************************************************
	    ATTENTION! Please answer the following quesiton in your lab report! Points will be allocated for the answers!
		 Hidden Question #1/2:
          What are the advantages and/or disadvantages of using a USB interface over PS/2 interface to
			 connect to the keyboard? List any two.  Give an answer in your Post-Lab.
     **************************************************************************************/
endmodule
